library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IM is
  port ( add  : in  STD_LOGIC_VECTOR(4 downto 0);
         instruction : out STD_LOGIC_VECTOR(31 downto 0));
end entity IM;

architecture dataflow of IM is
	 
    type mem_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
	 signal instrucmem : mem_array := (

	 "00000010011100101000100000100000", -- add $3, $2, $1
	 "00000010011100101000100000100010", -- sub $3, $2, $1
	 "00000010011100101000100000100101", -- or  $3, $2, $1
	 
	 "00000010001100101001100000100010", -- s
	 "00000100000000010000000001100100", 
	 "00000100000000100000000001100100", 
	 "00000000000000000000000000011001",
	 "00000000000000000000000000011000",
	 "00000000000000000000000000010111",
	 "00000000000000000000000000010110",
	 "00000000000000000000000000010101", -- 10
	 "00000000000000000000000000010100",
	 "00000000000000000000000000010011",
	 "00000000000000000000000000010010",
	 "00000000000000000000000000010001",
	 "00000000000000000000000000010000",
	 "00000000000000000000000000001111",
	 "00000000000000000000000000001110",
	 "00000000000000000000000000001101",
	 "00000000000000000000000000001100",
	 "00000000000000000000000000001011", -- 20
	 "00000000000000000000000000001010",
	 "00000000000000000000000000001001",
	 "00000000000000000000000000001000",
	 "00000000000000000000000000000111",
	 "00000000000000000000000000000110",
	 "00000000000000000000000000000101",
	 "00000000000000000000000000000100",
	 "00000000000000000000000000000011",  
	 "00000000000000000000000000000010",  
	 "00000000000000000000000000000001",  
	 "00000000000000000000000000000000"); 
BEGIN
    instruction <= instrucmem(TO_INTEGER(UNSIGNED(add)));
END dataflow;